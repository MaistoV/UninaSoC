`define TARGET_VIVADO
// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// Author: Florian Zaruba, ETH Zurich
// Date: 29.10.2018
// Description: Dummy circuit to mitigate Open Pin warnings

/* verilator lint_off UNUSED */
module unread (
    input logic d_i
);
    // Vivado treats this module as black box otherwise
`ifdef TARGET_VIVADO
    logic x;
    assign d_i = x;
`endif
endmodule
/* verilator lint_on UNUSED */